///////////////////////////
// WB Stage 
//////////////////////////
