//////////////////////////////////////////////////////
// Main CPU module                                 //
// This module will instantiate the other modules //
//                                               //
//////////////////////////////////////////////////
module CPU(
    .clk(clk),
    .rst_n(rst_n)
);
//We will need to instantiate wires between each pipeline
//stage and register instantiate the wires coming from each 
//stage or register in the specified section below

//IF Wires

//IF_ID_reg wires

//ID Wires

//ID_EX_reg wires

//EX_wires

//EX_MEM_reg wires

//MEM Wires

//MEM_WB_reg Wires

//WB Wires

//Hazard Unit Wires

//Forwarding Unit Wires

/////////////////////////////////
//Instantiate CPU Modules here//
///////////////////////////////
//IF Module

//IF_ID_reg Module

//ID Module

//ID_EX_reg Module

//EX Module

//EX_MEM_reg Module

//MEM Module

//MEM_WB_reg Module

//WB Module

//Hazard Unit 

//Forwarding Unit

endmodule
