//////////////////////////////////
// Module Name: MEM
// Author: Dustin R. Wiczek
// Module Summary: 
//
//////////////////////////////////
module MEM(
    input [31:0] mem_out,
    input




);


endmodule
//Line for revision controll version 1.0
